hviobj
